module top_module( output one );

// Insert your code here
    assign one = 1; //assign allows to drive an output continuously with a value, 十進位

endmodule
