module top_module(output zero);// Module body starts after semicolon
    //assign allows to drive an output continuously with a value
	assign zero = 0; //bits' decimal value
endmodule
