module top_module( input in, output out );
	assign out = in; // connect in to out
endmodule
